//------------------------------------------------------------------------
// Input Conditioner
//    1) Synchronizes input to clock domain
//    2) Debounces input
//    3) Creates pulses at edge transitions
//------------------------------------------------------------------------

module inputconditioner
(
input 	    clk,            // Clock domain to synchronize input to
input	    noisysignal,    // (Potentially) noisy input signal
output reg  conditioned = 0,    // Conditioned output signal
output reg  positiveedge = 0,   // 1 clk pulse at rising edge of conditioned
output reg  negativeedge = 0    // 1 clk pulse at falling edge of conditioned
);

/*Modify the module so that the positiveedge and negativeedge output signals
are correctly generated. These signals should be high for exactly one clock
period when conditioned has a positive/negative edge, starting in the same
clock period that conditioned transitions.

Note: There are several possible ways to generate the edge signals.
Remember that assign statements are continuous and operate on wires,
while assignments in always blocks (e.g. nonblocking <=) operate on regs.
*/

    parameter counterwidth = 3; // Counter size, in bits, >= log2(waittime)
    parameter waittime = 3;     // Debounce delay, in clock cycles

    reg[counterwidth-1:0] counter = 0;
    reg synchronizer0 = 0;
    reg synchronizer1 = 0;

    always @(posedge clk) begin
        positiveedge <= 0;
        negativeedge <= 0;
        if(conditioned == synchronizer1)
            counter <= 0;
        else begin
            if( counter == waittime) begin
                counter <= 0;
                conditioned <= synchronizer1;
                positiveedge <= synchronizer1;
                negativeedge <= !synchronizer1;
            end
            else
                counter <= counter+1;
        end
        synchronizer0 <= noisysignal;
        synchronizer1 <= synchronizer0;
    end
endmodule
