//------------------------------------------------------------------------
// Data Memory
//   Positive edge triggered
//   dataOut always has the value mem[address]
//   If writeEnable is true, writes dataIn to mem[address]
//------------------------------------------------------------------------

module finitestatemachine
(
    input  rising_sclk,
    input  conditioned_cs,
    input  shiftreg_out,
    output miso_bufe,
    output dm_we,
    output addr_we,
    output sr_we
);

    

endmodule
